
//-- Constants for obtaining standard BAURATES:
`define B115200 434
`define B57600 868
`define B38400 1302
`define B19200 2604
`define B9600 5208
`define B4800 10417
`define B2400 20833
`define B1200 41667
`define B600 83333
`define B300 166667